module backprop
  ();

   

endmodule: backprop
