module chip_interface;

    // uart_clock_divider -> goes to all next things
    // uart_recv
    // uart_protocol
    // control_unit

endmodule: chip_interface
