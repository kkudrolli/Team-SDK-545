module neuron
  (clk, rst, clear, );
   
   
endmodule: neuron
