module neuron
  (clk, rst_l, clear, );
   
   
endmodule: neuron
